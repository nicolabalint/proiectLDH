NAND3
.SUBCKT NAND3 1 2 3 7 6
MN1 6 1 5 0 CMOSN_35 L=0.35U W=1.32U
MN2 5 2 4 0 CMOSN_35 L=0.35U W=1.32U
MN3 4 3 0 0 CMOSN_35 L=0.35U W=1.32U
MP1 6 1 7 7 CMOSP_35 L=0.35U W=1.2U
MP2 6 2 7 7 CMOSP_35 L=0.35U W=1.2U
MP3 6 3 7 7 CMOSP_35 L=0.35U W=1.2U
.ENDS

VIN 1 0 0 PULSE(0 3.3 0 1N 1N 10N 20N)
VDD 10 0 3.3
X1 1 10 10 10 8 NAND3
CL 8 0 0.1P
.INC CMOS_035.txt

.TRAN 0.1N 20N 0 0.1N

.PROBE
.END