CIRCUIT
VD 14 0 0 PULSE(0 5V {TD} {TR} {TR} {PW1} 20n)
VCLK 16 0 0 PULSE(0 5V 2n {TR} {TR} {PW2} 10n)
VS 15 0 0 PULSE(0 5V 10N {TR} {TR} 100N 200N)
VDD 10 0 5

X1 14 20 19 10 21 INV3
X2 16 10 19 INV
X3 19 10 20 INV
X4 21 15 10 22 NAND2
X5 22 19 20  10 21 INV3
X6 22  19 20 10 23 INV3
X7 24 20 19 10 23 INV3
X8 23 15 10 24 NAND2
X9 24 10 25 INV
X10 24 10 18 INV
X11 25 10 17 INV

CL1 17 0 {CL}
CL2 18 0 {CL}

.inc "SUBCIRCUITE.txt"
.inc "CMOS_HP_05_T49G.txt"
.PARAM CL=0.1p
.PARAM TR=50p
.PARAM TD=0
.PARAM PW1=10N
.PARAM PW2=5N
*.STEP PARAM TD 0 10N 0.1N
*.STEP PARAM PW1 6.99N 7N 0.001N
.STEP PARAM PW2 0.2n 0.25n 0.001n
.tran 0.1n 60n
.probe
.end
