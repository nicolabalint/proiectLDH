NOR3
.SUBCKT NOR3 1 2 3 7 4
MN1 4 1 0 0 CMOSN_35 L=0.35U W=0.8U
MN2 4 2 0 0 CMOSN_35 L=0.35U W=0.8U
MN3 4 3 0 0 CMOSN_35 L=0.35U W=0.8U
MP1 6 1 7 7 CMOSP_35 L=0.35U W=6.48U
MP2 5 2 6 7 CMOSP_35 L=0.35U W=6.48U
MP3 4 3 5 7 CMOSP_35 L=0.35U W=6.48U
.ENDS

VIN 1 0 0 PULSE(0 3.3 0 1N 1N 10N 20N)
VDD 10 0 3.3
X1 1 0 0 10 8 NOR3
CL 8 0 0.1P
.INC CMOS_035.txt

.TRAN 0.1N 20N 0 0.1N

.PROBE
.END